
module pll (
	);	

endmodule
