	component pll is
	end component pll;

	u0 : component pll
		port map (
		);

